LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY fcoc IS 
	PORT (A1,B1,S0:IN STD_LOGIC;
				Y1:OUT STD_LOGIC);
END ENTITY fcoc;
ARCHITECTURE BHV OF fcoc IS
	BEGIN
	
END ARCHITECTURE BHV;